//`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////////
//// Company: 
//// Engineer: 
//// 
//// Create Date: 09.10.2024 21:25:14
//// Design Name: 
//// Module Name: mixColumnstb
//// Project Name: 
//// Target Devices: 
//// Tool Versions: 
//// Description: 
//// 
//// Dependencies: 
//// 
//// Revision:
//// Revision 0.01 - File Created
//// Additional Comments:
//// 
////////////////////////////////////////////////////////////////////////////////////


//module mixColumns_tb;
//    reg [7:0] state [0:3][0:3];
//    wire [7:0] out [0:3][0:3];
    
//    mixColumns dut (
//        .state(state),
//        .out(out)
//    );

//    initial begin
//        state[0][0] = 8'h63; state[0][1] = 8'hA5; state[0][2] = 8'hC3; state[0][3] = 8'hFD;
//        state[1][0] = 8'h8F; state[1][1] = 8'h71; state[1][2] = 8'h04; state[1][3] = 8'h27;
//        state[2][0] = 8'h18; state[2][1] = 8'h26; state[2][2] = 8'h63; state[2][3] = 8'hFE;
//        state[3][0] = 8'h34; state[3][1] = 8'h37; state[3][2] = 8'h61; state[3][3] = 8'h0A;
//        #10;
//        $finish;
//    end
//endmodule

