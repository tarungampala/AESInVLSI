//`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////////
//// Company: 
//// Engineer: 
//// 
//// Create Date: 09.10.2024 19:49:08
//// Design Name: 
//// Module Name: shiftrowstb
//// Project Name: 
//// Target Devices: 
//// Tool Versions: 
//// Description: 
//// 
//// Dependencies: 
//// 
//// Revision:
//// Revision 0.01 - File Created
//// Additional Comments:
//// 
////////////////////////////////////////////////////////////////////////////////////


//module shiftrowstb();
//    reg [7:0] in [0:3][0:3];
//    wire [7:0] out [0:3][0:3];
    
//    shiftRows dut (.in(in), .out(out));
    
//    initial begin
//        in[0][0] = 8'h63; in[0][1] = 8'hA5; in[0][2] = 8'hC3; in[0][3] = 8'hFD;
//        in[1][0] = 8'h27; in[1][1] = 8'h8F; in[1][2] = 8'h71; in[1][3] = 8'h04;
//        in[2][0] = 8'h63; in[2][1] = 8'hFE; in[2][2] = 8'h18; in[2][3] = 8'h26;
//        in[3][0] = 8'h37; in[3][1] = 8'h61; in[3][2] = 8'h0A; in[3][3] = 8'h34;
        
//        #5;
//        $finish();
//    end
    
//endmodule
