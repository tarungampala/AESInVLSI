//`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////////
//// Company: 
//// Engineer: 
//// 
//// Create Date: 09.10.2024 18:59:23
//// Design Name: 
//// Module Name: roundkeytb
//// Project Name: 
//// Target Devices: 
//// Tool Versions: 
//// Description: 
//// 
//// Dependencies: 
//// 
//// Revision:
//// Revision 0.01 - File Created
//// Additional Comments:
//// 
////////////////////////////////////////////////////////////////////////////////////


//module roundkeytb();
//    reg [0:7] in [0:3][0:3];
//    reg [0:7] key [0:3][0:3];
//    wire [0:7] out [0:3][0:3];
    
//    roundkey dut (.in(in), .key(key), .out(out));
    
//    initial begin
//        in[0][0] = 8'h54; in[0][1] = 8'h41; in[0][2] = 8'h52; in[0][3] = 8'h55;
//        in[1][0] = 8'h4E; in[1][1] = 8'h53; in[1][2] = 8'h41; in[1][3] = 8'h49;
//        in[2][0] = 8'h20; in[2][1] = 8'h47; in[2][2] = 8'h41; in[2][3] = 8'h4D;
//        in[3][0] = 8'h50; in[3][1] = 8'h41; in[3][2] = 8'h4C; in[3][3] = 8'h41;
       
//        key[0][0] = 8'h54; key[0][1] = 8'h68; key[0][2] = 8'h61; key[0][3] = 8'h74;
//        key[1][0] = 8'h73; key[1][1] = 8'h20; key[1][2] = 8'h6D; key[1][3] = 8'h79;
//        key[2][0] = 8'h20; key[2][1] = 8'h4B; key[2][2] = 8'h75; key[2][3] = 8'h6E;
//        key[3][0] = 8'h67; key[3][1] = 8'h20; key[3][2] = 8'h46; key[3][3] = 8'h75; 
        
//        #5;
//        $finish();
//    end
//endmodule
