//`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////////
//// Company: 
//// Engineer: 
//// 
//// Create Date: 09.10.2024 20:09:33
//// Design Name: 
//// Module Name: subBytestb
//// Project Name: 
//// Target Devices: 
//// Tool Versions: 
//// Description: 
//// 
//// Dependencies: 
//// 
//// Revision:
//// Revision 0.01 - File Created
//// Additional Comments:
//// 
////////////////////////////////////////////////////////////////////////////////////


//module subBytestb();
//    logic [7:0] state [0:3][0:3];
//    logic [7:0] outState [0:3][0:3];

//    // Instantiate the SubBytes module
//    subBytes dut (.state(state), .outState(outState));

//    initial begin
//        state[0][0] = 8'h00;
//        state[0][1] = 8'h29;
//        state[0][2] = 8'h33;
//        state[0][3] = 8'h21;
        
//        state[1][0] = 8'h3D;
//        state[1][1] = 8'h73;
//        state[1][2] = 8'h2C;
//        state[1][3] = 8'h30;
        
//        state[2][0] = 8'h00;
//        state[2][1] = 8'h0C;
//        state[2][2] = 8'h34;
//        state[2][3] = 8'h23;
        
//        state[3][0] = 8'h37;
//        state[3][1] = 8'h61;
//        state[3][2] = 8'h0A;
//        state[3][3] = 8'h34;

//        #1;
//        $finish();
//   end
//endmodule
